module runtime

fn current_process_mem_usage_mac() u32 {
	return 0
}